-- VJTAG.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity VJTAG is
	port (
		tdi                : out std_logic;                                       -- jtag.tdi
		tdo                : in  std_logic                    := '0';             --     .tdo
		ir_in              : out std_logic_vector(0 downto 0);                    --     .ir_in
		ir_out             : in  std_logic_vector(0 downto 0) := (others => '0'); --     .ir_out
		virtual_state_cdr  : out std_logic;                                       --     .virtual_state_cdr
		virtual_state_sdr  : out std_logic;                                       --     .virtual_state_sdr
		virtual_state_e1dr : out std_logic;                                       --     .virtual_state_e1dr
		virtual_state_pdr  : out std_logic;                                       --     .virtual_state_pdr
		virtual_state_e2dr : out std_logic;                                       --     .virtual_state_e2dr
		virtual_state_udr  : out std_logic;                                       --     .virtual_state_udr
		virtual_state_cir  : out std_logic;                                       --     .virtual_state_cir
		virtual_state_uir  : out std_logic;                                       --     .virtual_state_uir
		tms                : out std_logic;                                       --     .tms
		jtag_state_tlr     : out std_logic;                                       --     .jtag_state_tlr
		jtag_state_rti     : out std_logic;                                       --     .jtag_state_rti
		jtag_state_sdrs    : out std_logic;                                       --     .jtag_state_sdrs
		jtag_state_cdr     : out std_logic;                                       --     .jtag_state_cdr
		jtag_state_sdr     : out std_logic;                                       --     .jtag_state_sdr
		jtag_state_e1dr    : out std_logic;                                       --     .jtag_state_e1dr
		jtag_state_pdr     : out std_logic;                                       --     .jtag_state_pdr
		jtag_state_e2dr    : out std_logic;                                       --     .jtag_state_e2dr
		jtag_state_udr     : out std_logic;                                       --     .jtag_state_udr
		jtag_state_sirs    : out std_logic;                                       --     .jtag_state_sirs
		jtag_state_cir     : out std_logic;                                       --     .jtag_state_cir
		jtag_state_sir     : out std_logic;                                       --     .jtag_state_sir
		jtag_state_e1ir    : out std_logic;                                       --     .jtag_state_e1ir
		jtag_state_pir     : out std_logic;                                       --     .jtag_state_pir
		jtag_state_e2ir    : out std_logic;                                       --     .jtag_state_e2ir
		jtag_state_uir     : out std_logic;                                       --     .jtag_state_uir
		tck                : out std_logic                                        --  tck.clk
	);
end entity VJTAG;

architecture rtl of VJTAG is
	component sld_virtual_jtag is
		generic (
			sld_auto_instance_index : string  := "YES";
			sld_instance_index      : integer := 0;
			sld_ir_width            : integer := 1
		);
		port (
			tdi                : out std_logic;                                       -- tdi
			tdo                : in  std_logic                    := 'X';             -- tdo
			ir_in              : out std_logic_vector(0 downto 0);                    -- ir_in
			ir_out             : in  std_logic_vector(0 downto 0) := (others => 'X'); -- ir_out
			virtual_state_cdr  : out std_logic;                                       -- virtual_state_cdr
			virtual_state_sdr  : out std_logic;                                       -- virtual_state_sdr
			virtual_state_e1dr : out std_logic;                                       -- virtual_state_e1dr
			virtual_state_pdr  : out std_logic;                                       -- virtual_state_pdr
			virtual_state_e2dr : out std_logic;                                       -- virtual_state_e2dr
			virtual_state_udr  : out std_logic;                                       -- virtual_state_udr
			virtual_state_cir  : out std_logic;                                       -- virtual_state_cir
			virtual_state_uir  : out std_logic;                                       -- virtual_state_uir
			tms                : out std_logic;                                       -- tms
			jtag_state_tlr     : out std_logic;                                       -- jtag_state_tlr
			jtag_state_rti     : out std_logic;                                       -- jtag_state_rti
			jtag_state_sdrs    : out std_logic;                                       -- jtag_state_sdrs
			jtag_state_cdr     : out std_logic;                                       -- jtag_state_cdr
			jtag_state_sdr     : out std_logic;                                       -- jtag_state_sdr
			jtag_state_e1dr    : out std_logic;                                       -- jtag_state_e1dr
			jtag_state_pdr     : out std_logic;                                       -- jtag_state_pdr
			jtag_state_e2dr    : out std_logic;                                       -- jtag_state_e2dr
			jtag_state_udr     : out std_logic;                                       -- jtag_state_udr
			jtag_state_sirs    : out std_logic;                                       -- jtag_state_sirs
			jtag_state_cir     : out std_logic;                                       -- jtag_state_cir
			jtag_state_sir     : out std_logic;                                       -- jtag_state_sir
			jtag_state_e1ir    : out std_logic;                                       -- jtag_state_e1ir
			jtag_state_pir     : out std_logic;                                       -- jtag_state_pir
			jtag_state_e2ir    : out std_logic;                                       -- jtag_state_e2ir
			jtag_state_uir     : out std_logic;                                       -- jtag_state_uir
			tck                : out std_logic                                        -- clk
		);
	end component sld_virtual_jtag;

begin

	virtual_jtag_0 : component sld_virtual_jtag
		generic map (
			sld_auto_instance_index => "YES",
			sld_instance_index      => 0,
			sld_ir_width            => 1
		)
		port map (
			tdi                => tdi,                -- jtag.tdi
			tdo                => tdo,                --     .tdo
			ir_in              => ir_in,              --     .ir_in
			ir_out             => ir_out,             --     .ir_out
			virtual_state_cdr  => virtual_state_cdr,  --     .virtual_state_cdr
			virtual_state_sdr  => virtual_state_sdr,  --     .virtual_state_sdr
			virtual_state_e1dr => virtual_state_e1dr, --     .virtual_state_e1dr
			virtual_state_pdr  => virtual_state_pdr,  --     .virtual_state_pdr
			virtual_state_e2dr => virtual_state_e2dr, --     .virtual_state_e2dr
			virtual_state_udr  => virtual_state_udr,  --     .virtual_state_udr
			virtual_state_cir  => virtual_state_cir,  --     .virtual_state_cir
			virtual_state_uir  => virtual_state_uir,  --     .virtual_state_uir
			tms                => tms,                --     .tms
			jtag_state_tlr     => jtag_state_tlr,     --     .jtag_state_tlr
			jtag_state_rti     => jtag_state_rti,     --     .jtag_state_rti
			jtag_state_sdrs    => jtag_state_sdrs,    --     .jtag_state_sdrs
			jtag_state_cdr     => jtag_state_cdr,     --     .jtag_state_cdr
			jtag_state_sdr     => jtag_state_sdr,     --     .jtag_state_sdr
			jtag_state_e1dr    => jtag_state_e1dr,    --     .jtag_state_e1dr
			jtag_state_pdr     => jtag_state_pdr,     --     .jtag_state_pdr
			jtag_state_e2dr    => jtag_state_e2dr,    --     .jtag_state_e2dr
			jtag_state_udr     => jtag_state_udr,     --     .jtag_state_udr
			jtag_state_sirs    => jtag_state_sirs,    --     .jtag_state_sirs
			jtag_state_cir     => jtag_state_cir,     --     .jtag_state_cir
			jtag_state_sir     => jtag_state_sir,     --     .jtag_state_sir
			jtag_state_e1ir    => jtag_state_e1ir,    --     .jtag_state_e1ir
			jtag_state_pir     => jtag_state_pir,     --     .jtag_state_pir
			jtag_state_e2ir    => jtag_state_e2ir,    --     .jtag_state_e2ir
			jtag_state_uir     => jtag_state_uir,     --     .jtag_state_uir
			tck                => tck                 --  tck.clk
		);

end architecture rtl; -- of VJTAG
